package test_order_pkg is

  constant THE_TRUTH : integer := 42;

end package test_order_pkg;
